version https://git-lfs.github.com/spec/v1
oid sha256:059e6ceb1b7d88363a654934bbcb258845923cb936c1f2370b5b861244504b5f
size 11803
