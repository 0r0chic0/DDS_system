version https://git-lfs.github.com/spec/v1
oid sha256:a7649b25a40bd13fbbff2a94ee9030e017c4c3f22ef4c9d46192a78e308d74b3
size 1598
