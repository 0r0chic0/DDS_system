version https://git-lfs.github.com/spec/v1
oid sha256:976b292f813aae949e894517da1d0085d5cb31d6de74619b5bfd41417e4acecd
size 10715
