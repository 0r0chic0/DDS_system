version https://git-lfs.github.com/spec/v1
oid sha256:b4bcced5fc46d3d83ad2da086fa461f9179db92f6b5fbd78695db0d472e9430c
size 26475
