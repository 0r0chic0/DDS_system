version https://git-lfs.github.com/spec/v1
oid sha256:3904c8d8e59375aadce1c76e99214c7af158bf65eb0a09535580077397fcf7c6
size 3450
