version https://git-lfs.github.com/spec/v1
oid sha256:4aef61d2ff28cb78abfd965212a679857aeef796ca8f6bf8ae9bd5c9d7cf98da
size 3780
