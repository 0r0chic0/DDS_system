version https://git-lfs.github.com/spec/v1
oid sha256:2955b11424ff31cc94f15d40ee86153603ed158842c4e3b788599e628ee99565
size 7914
