version https://git-lfs.github.com/spec/v1
oid sha256:60b1f8f15371a2b069fd708cf2e8929ba11289a0f7fb45d6d8108c03eb6a192b
size 15339
