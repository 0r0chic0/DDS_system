version https://git-lfs.github.com/spec/v1
oid sha256:45a5b9f8217fbe53b67c11e8174f8e3c71dc1f1219f7774b2f61c63292b1a43c
size 8224
