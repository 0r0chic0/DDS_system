version https://git-lfs.github.com/spec/v1
oid sha256:eb421650a9b0011f54451e1b97d167bd57fb0a3ea97c82c50a2a1a118430cd82
size 4700
