version https://git-lfs.github.com/spec/v1
oid sha256:ab455bb0dbed5d22a69f7b1735a19a0a3bf4229b894c3a41e6dca2e2f4a6e541
size 7718
