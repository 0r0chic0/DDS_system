version https://git-lfs.github.com/spec/v1
oid sha256:b908b871447072c9c216ae742601e0e7a9677b2b32a90233ef8865b4f67013a8
size 3458
