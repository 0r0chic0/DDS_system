version https://git-lfs.github.com/spec/v1
oid sha256:387ab4a6f2aef1562650286364bbf09ad1c989583bb0d7bdb36395338866dc5e
size 8006
