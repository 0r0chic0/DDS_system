version https://git-lfs.github.com/spec/v1
oid sha256:f0a01ef6db58433f6265e95d5f081db4c326db6a9d0d779c52fac63bad6be0d5
size 29775
