version https://git-lfs.github.com/spec/v1
oid sha256:edbcbb65be4970ed4c4b312d0b60d3f1ef859daccdeaf19c016b66175b704c36
size 3715
