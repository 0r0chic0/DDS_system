version https://git-lfs.github.com/spec/v1
oid sha256:0db28d28d6727187fc30c33c6299e01cb60b1d78804869d116eb401588bad75c
size 11051
