version https://git-lfs.github.com/spec/v1
oid sha256:0444d5db7c42b61b6d0df0e52c41e64c126e07eec1cbd6239f48d5c6bb39c2d5
size 3458
