version https://git-lfs.github.com/spec/v1
oid sha256:31b4bdbe593430fdac412f39aeed501284d5d1c759ec41dc743ba4ce8b51a2cf
size 3772
