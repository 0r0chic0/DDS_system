version https://git-lfs.github.com/spec/v1
oid sha256:e559175d82016554f9589fd9dc1118e2b8583bfbefb8269f8d0a3da9be32ee99
size 7908
