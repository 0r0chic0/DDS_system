version https://git-lfs.github.com/spec/v1
oid sha256:6583ce871291d5d576bea16d0af9d280ee0ac077fbafed22c516f654846eb0e8
size 3718
