version https://git-lfs.github.com/spec/v1
oid sha256:c4adc73995105c99c5ff653fab5a0014bd60caec91ccf21b18ca077996393b9a
size 7546
