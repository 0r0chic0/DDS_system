version https://git-lfs.github.com/spec/v1
oid sha256:ad52a29d0dae57e27da658b28f7cb40c8eeab3208656b818fc972876cdb7dab2
size 4079
