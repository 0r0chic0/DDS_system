version https://git-lfs.github.com/spec/v1
oid sha256:2691b77d7c9e91a954eabad93a5c9d027c5793aa8ff1153574d1e8ccf519aaad
size 43369
