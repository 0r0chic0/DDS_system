version https://git-lfs.github.com/spec/v1
oid sha256:9cf36ef68b2c2ec1ba540d336480ce2c409375df7c94fa4df1fbcc3ec55fdaf5
size 2012
