version https://git-lfs.github.com/spec/v1
oid sha256:6fadf564af80ba4350c9962cf970376298afbcd18f867945372783d2bb077581
size 11773
