version https://git-lfs.github.com/spec/v1
oid sha256:b050445b50f768d4617672926f124e64e86df05c8e57eed1c59b985f0a8bc145
size 3458
