version https://git-lfs.github.com/spec/v1
oid sha256:dc184070c154d7db744490e7581a1da3c9918965dfef5596772695b579bd6fed
size 18530
